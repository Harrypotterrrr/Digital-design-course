`timescale 1ns / 1ps
module pcreg(
    input clk, //1 λ���룬�Ĵ���ʱ���źţ�������ʱΪ PC �Ĵ�����ֵ
    input rst, //1 λ���룬 �첽�����źţ��ߵ�ƽʱ�� PC �Ĵ�������
    //ע���� ena �ź���Чʱ�� rst Ҳ�������üĴ���
    input ena, //1 λ����,��Ч�źŸߵ�ƽʱ PC �Ĵ������� data_in
    //��ֵ�����򱣳�ԭ�����
    input [31:0] data_in, //32 λ���룬�������ݽ�������Ĵ����ڲ�
    output wire [31:0] data_out //32 λ���������ʱʼ����� PC
    //�Ĵ����ڲ��洢��ֵ
);
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test0(
            .CLK(clk),
            .D(data_in[0]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[0])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test1(
            .CLK(clk),
            .D(data_in[1]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[1])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test2(
            .CLK(clk),
            .D(data_in[2]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[2])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test3(
            .CLK(clk),
            .D(data_in[3]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[3])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test4(
            .CLK(clk),
            .D(data_in[4]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[4])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test5(
            .CLK(clk),
            .D(data_in[5]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[5])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test6(
            .CLK(clk),
            .D(data_in[6]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[6])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test7(
            .CLK(clk),
            .D(data_in[7]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[7])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test8(
            .CLK(clk),
            .D(data_in[8]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[8])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test9(
            .CLK(clk),
            .D(data_in[9]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[9])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test10(
            .CLK(clk),
            .D(data_in[10]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[10])
        );
        Asynchronous_D_pcreg      
        Asynchronous_D_pcreg_test11(
            .CLK(clk),
            .D(data_in[11]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[11])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test12(
            .CLK(clk),
            .D(data_in[12]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[12])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test13(
            .CLK(clk),
            .D(data_in[13]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[13])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test14(
            .CLK(clk),
            .D(data_in[14]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[14])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test15(
            .CLK(clk),
            .D(data_in[15]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[15])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test16(
            .CLK(clk),
            .D(data_in[16]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[16])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test17(
            .CLK(clk),
            .D(data_in[17]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[17])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test18(
            .CLK(clk),
            .D(data_in[18]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[18])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test19(
            .CLK(clk),
            .D(data_in[19]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[19])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test20(
            .CLK(clk),
            .D(data_in[20]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[20])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test21(
            .CLK(clk),
            .D(data_in[21]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[21])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test22(
            .CLK(clk),
            .D(data_in[22]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[22])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test23(
            .CLK(clk),
            .D(data_in[23]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[23])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test24(
            .CLK(clk),
            .D(data_in[24]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[24])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test25(
            .CLK(clk),
            .D(data_in[25]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[25])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test26(
            .CLK(clk),
            .D(data_in[26]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[26])
        );
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test27(
            .CLK(clk),
            .D(data_in[27]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[27])
        );
        Asynchronous_D_pcreg      
        Asynchronous_D_pcreg_test28(
            .CLK(clk),
            .D(data_in[28]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[28])
        );   
        Asynchronous_D_pcreg   
        Asynchronous_D_pcreg_test29(
            .CLK(clk),
            .D(data_in[29]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[29])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test30(
            .CLK(clk),
            .D(data_in[30]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[30])
        );      
        Asynchronous_D_pcreg
        Asynchronous_D_pcreg_test31(
            .CLK(clk),
            .D(data_in[31]),
            .RST_n(rst),
            .ena(ena),
            .Out(data_out[31])
        );      

endmodule
